module ram_1KB_instruction #(  parameter MEM_FILE   = "")
(i_clk, i_rst, i_address, o_data);

input logic i_clk;
input logic i_rst;
//input logic i_wren;
input logic [7:0] i_address;
//input logic [31:0] i_data;
output logic [31:0] o_data;
logic [31:0] mem [0:255]; 


    initial begin
        if (MEM_FILE != "") begin
            $readmemh(MEM_FILE, mem);
        end
    end

always_ff @(posedge i_clk or negedge i_rst) begin
    if (!i_rst) begin
        mem[0] <= 32'b0;
        mem[1] <= 32'b0;
        mem[2] <= 32'b0;
        mem[3] <= 32'b0;
        mem[4] <= 32'b0;
        mem[5] <= 32'b0;
        mem[6] <= 32'b0;
        mem[7] <= 32'b0;
        mem[8] <= 32'b0;
        mem[9] <= 32'b0;
        mem[10] <= 32'b0;
        mem[11] <= 32'b0;
        mem[12] <= 32'b0;
        mem[13] <= 32'b0;
        mem[14] <= 32'b0;
        mem[15] <= 32'b0;
        mem[16] <= 32'b0;
        mem[17] <= 32'b0;
        mem[18] <= 32'b0;
        mem[19] <= 32'b0;
        mem[20] <= 32'b0;
        mem[21] <= 32'b0;
        mem[22] <= 32'b0;
        mem[23] <= 32'b0;
        mem[24] <= 32'b0;
        mem[25] <= 32'b0;
        mem[26] <= 32'b0;
        mem[27] <= 32'b0;
        mem[28] <= 32'b0;
        mem[29] <= 32'b0;
        mem[30] <= 32'b0;
        mem[31] <= 32'b0;
        mem[32] <= 32'b0;
        mem[33] <= 32'b0;
        mem[34] <= 32'b0;
        mem[35] <= 32'b0;
        mem[36] <= 32'b0;
        mem[37] <= 32'b0;
        mem[38] <= 32'b0;
        mem[39] <= 32'b0;
        mem[40] <= 32'b0;
        mem[41] <= 32'b0;
        mem[42] <= 32'b0;
        mem[43] <= 32'b0;
        mem[44] <= 32'b0;
        mem[45] <= 32'b0;
        mem[46] <= 32'b0;
        mem[47] <= 32'b0;
        mem[48] <= 32'b0;
        mem[49] <= 32'b0;
        mem[50] <= 32'b0;
        mem[51] <= 32'b0;
        mem[52] <= 32'b0;
        mem[53] <= 32'b0;
        mem[54] <= 32'b0;
        mem[55] <= 32'b0;
        mem[56] <= 32'b0;
        mem[57] <= 32'b0;
        mem[58] <= 32'b0;
        mem[59] <= 32'b0;
        mem[60] <= 32'b0;
        mem[61] <= 32'b0;
        mem[62] <= 32'b0;
        mem[63] <= 32'b0;
        mem[64] <= 32'b0;
        mem[65] <= 32'b0;
        mem[66] <= 32'b0;
        mem[67] <= 32'b0;
        mem[68] <= 32'b0;
        mem[69] <= 32'b0;
        mem[70] <= 32'b0;
        mem[71] <= 32'b0;
        mem[72] <= 32'b0;
        mem[73] <= 32'b0;
        mem[74] <= 32'b0;
        mem[75] <= 32'b0;
        mem[76] <= 32'b0;
        mem[77] <= 32'b0;
        mem[78] <= 32'b0;
        mem[79] <= 32'b0;
        mem[80] <= 32'b0;
        mem[81] <= 32'b0;
        mem[82] <= 32'b0;
        mem[83] <= 32'b0;
        mem[84] <= 32'b0;
        mem[85] <= 32'b0;
        mem[86] <= 32'b0;
        mem[87] <= 32'b0;
        mem[88] <= 32'b0;
        mem[89] <= 32'b0;
        mem[90] <= 32'b0;
        mem[91] <= 32'b0;
        mem[92] <= 32'b0;
        mem[93] <= 32'b0;
        mem[94] <= 32'b0;
        mem[95] <= 32'b0;
        mem[96] <= 32'b0;
        mem[97] <= 32'b0;
        mem[98] <= 32'b0;
        mem[99] <= 32'b0;
        mem[100] <= 32'b0;
        mem[101] <= 32'b0;
        mem[102] <= 32'b0;
        mem[103] <= 32'b0;
        mem[104] <= 32'b0;
        mem[105] <= 32'b0;
        mem[106] <= 32'b0;
        mem[107] <= 32'b0;
        mem[108] <= 32'b0;
        mem[109] <= 32'b0;
        mem[110] <= 32'b0;
        mem[111] <= 32'b0;
        mem[112] <= 32'b0;
        mem[113] <= 32'b0;
        mem[114] <= 32'b0;
        mem[115] <= 32'b0;
        mem[116] <= 32'b0;
        mem[117] <= 32'b0;
        mem[118] <= 32'b0;
        mem[119] <= 32'b0;
        mem[120] <= 32'b0;
        mem[121] <= 32'b0;
        mem[122] <= 32'b0;
        mem[123] <= 32'b0;
        mem[124] <= 32'b0;
        mem[125] <= 32'b0;
        mem[126] <= 32'b0;
        mem[127] <= 32'b0;
        mem[128] <= 32'b0;
        mem[129] <= 32'b0;
        mem[130] <= 32'b0;
        mem[131] <= 32'b0;
        mem[132] <= 32'b0;
        mem[133] <= 32'b0;
        mem[134] <= 32'b0;
        mem[135] <= 32'b0;
        mem[136] <= 32'b0;
        mem[137] <= 32'b0;
        mem[138] <= 32'b0;
        mem[139] <= 32'b0;
        mem[140] <= 32'b0;
        mem[141] <= 32'b0;
        mem[142] <= 32'b0;
        mem[143] <= 32'b0;
        mem[144] <= 32'b0;
        mem[145] <= 32'b0;
        mem[146] <= 32'b0;
        mem[147] <= 32'b0;
        mem[148] <= 32'b0;
        mem[149] <= 32'b0;
        mem[150] <= 32'b0;
        mem[151] <= 32'b0;
        mem[152] <= 32'b0;
        mem[153] <= 32'b0;
        mem[154] <= 32'b0;
        mem[155] <= 32'b0;
        mem[156] <= 32'b0;
        mem[157] <= 32'b0;
        mem[158] <= 32'b0;
        mem[159] <= 32'b0;
        mem[160] <= 32'b0;
        mem[161] <= 32'b0;
        mem[162] <= 32'b0;
        mem[163] <= 32'b0;
        mem[164] <= 32'b0;
        mem[165] <= 32'b0;
        mem[166] <= 32'b0;
        mem[167] <= 32'b0;
        mem[168] <= 32'b0;
        mem[169] <= 32'b0;
        mem[170] <= 32'b0;
        mem[171] <= 32'b0;
        mem[172] <= 32'b0;
        mem[173] <= 32'b0;
        mem[174] <= 32'b0;
        mem[175] <= 32'b0;
        mem[176] <= 32'b0;
        mem[177] <= 32'b0;
        mem[178] <= 32'b0;
        mem[179] <= 32'b0;
        mem[180] <= 32'b0;
        mem[181] <= 32'b0;
        mem[182] <= 32'b0;
        mem[183] <= 32'b0;
        mem[184] <= 32'b0;
        mem[185] <= 32'b0;
        mem[186] <= 32'b0;
        mem[187] <= 32'b0;
        mem[188] <= 32'b0;
        mem[189] <= 32'b0;
        mem[190] <= 32'b0;
        mem[191] <= 32'b0;
        mem[192] <= 32'b0;
        mem[193] <= 32'b0;
        mem[194] <= 32'b0;
        mem[195] <= 32'b0;
        mem[196] <= 32'b0;
        mem[197] <= 32'b0;
        mem[198] <= 32'b0;
        mem[199] <= 32'b0;
        mem[200] <= 32'b0;
        mem[201] <= 32'b0;
        mem[202] <= 32'b0;
        mem[203] <= 32'b0;
        mem[204] <= 32'b0;
        mem[205] <= 32'b0;
        mem[206] <= 32'b0;
        mem[207] <= 32'b0;
        mem[208] <= 32'b0;
        mem[209] <= 32'b0;
        mem[210] <= 32'b0;
        mem[211] <= 32'b0;
        mem[212] <= 32'b0;
        mem[213] <= 32'b0;
        mem[214] <= 32'b0;
        mem[215] <= 32'b0;
        mem[216] <= 32'b0;
        mem[217] <= 32'b0;
        mem[218] <= 32'b0;
        mem[219] <= 32'b0;
        mem[220] <= 32'b0;
        mem[221] <= 32'b0;
        mem[222] <= 32'b0;
        mem[223] <= 32'b0;
        mem[224] <= 32'b0;
        mem[225] <= 32'b0;
        mem[226] <= 32'b0;
        mem[227] <= 32'b0;
        mem[228] <= 32'b0;
        mem[229] <= 32'b0;
        mem[230] <= 32'b0;
        mem[231] <= 32'b0;
        mem[232] <= 32'b0;
        mem[233] <= 32'b0;
        mem[234] <= 32'b0;
        mem[235] <= 32'b0;
        mem[236] <= 32'b0;
        mem[237] <= 32'b0;
        mem[238] <= 32'b0;
        mem[239] <= 32'b0;
        mem[240] <= 32'b0;
        mem[241] <= 32'b0;
        mem[242] <= 32'b0;
        mem[243] <= 32'b0;
        mem[244] <= 32'b0;
        mem[245] <= 32'b0;
        mem[246] <= 32'b0;
        mem[247] <= 32'b0;
        mem[248] <= 32'b0;
        mem[249] <= 32'b0;
        mem[250] <= 32'b0;
        mem[251] <= 32'b0;
        mem[252] <= 32'b0;
        mem[253] <= 32'b0;
        mem[254] <= 32'b0;
        mem[255] <= 32'b0;
    end /*else if (i_wren) begin
        mem[i_address] <= i_data;
    end */
end 

always_comb begin
    o_data = mem[i_address];
end


endmodule         